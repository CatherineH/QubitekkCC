// megafunction wizard: %LPM_MUX%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: chan_mux.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.1.0 Build 162 10/23/2013 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module chan_mux (
	data0x,
	data1x,
	data2x,
	sel,
	result);

	input	[21:0]  data0x;
	input	[21:0]  data1x;
	input	[21:0]  data2x;
	input	[1:0]  sel;
	output	[21:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "3"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "22"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "2"
// Retrieval info: USED_PORT: data0x 0 0 22 0 INPUT NODEFVAL "data0x[21..0]"
// Retrieval info: USED_PORT: data1x 0 0 22 0 INPUT NODEFVAL "data1x[21..0]"
// Retrieval info: USED_PORT: data2x 0 0 22 0 INPUT NODEFVAL "data2x[21..0]"
// Retrieval info: USED_PORT: result 0 0 22 0 OUTPUT NODEFVAL "result[21..0]"
// Retrieval info: USED_PORT: sel 0 0 2 0 INPUT NODEFVAL "sel[1..0]"
// Retrieval info: CONNECT: @data 0 0 22 0 data0x 0 0 22 0
// Retrieval info: CONNECT: @data 0 0 22 22 data1x 0 0 22 0
// Retrieval info: CONNECT: @data 0 0 22 44 data2x 0 0 22 0
// Retrieval info: CONNECT: @sel 0 0 2 0 sel 0 0 2 0
// Retrieval info: CONNECT: result 0 0 22 0 @result 0 0 22 0
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL chan_mux_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
